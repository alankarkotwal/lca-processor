`ifndef _PIPELINE_REGS
`define _PIPELINE_REGS

module pipeline_reg1(); // First pipeline register

endmodule


module pipeline_reg2();

endmodule


module pipeline_reg3();

endmodule


module pipeline_reg4();

endmodule


module pipeline_reg5();

endmodule

`endif
