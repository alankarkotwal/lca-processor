`ifndef _REG_READ
`define _REG_READ

module reg_read();

endmodule

`endif
