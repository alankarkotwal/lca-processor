`ifndef _EXECUTE
`define _EXECUTE

module execute();

	

endmodule

`endif
