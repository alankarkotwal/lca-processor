`ifndef _LCA_PROCESSOR
`define _LCA_PROCESSOR

`include "../pipeline/pipeline_regs.v"
`include "../pipeline/fetch.v"

module lca_processor();

endmodule

`endif
