`ifndef _MEM_ACCESS
`define _MEM_ACCESS

module mem_access();

	

endmodule

`endif
