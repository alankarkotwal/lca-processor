`ifndef _LCA_PROCESSOR
`define _LCA_PROCESSOR

module lca_processor();

endmodule

`endif
