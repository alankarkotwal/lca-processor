`ifndef _DECODE
`define _DECODE

module decode();

endmodule

`endif
