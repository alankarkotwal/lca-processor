`ifndef _WRITE_BACK
`define _WRITE_BACK

module write_back();

endmodule

`endif
